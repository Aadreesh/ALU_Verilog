`include "or.v"
module or_all
{
    input [31:0] a, b,
    output [31:0] out
};
    or d0(y[0],a[0],b[0]);
    or d1(y[1],a[1],b[1]);
    or d2(y[2],a[2],b[2]);
    or d3(y[3],a[3],b[3]);
    or d4(y[4],a[4],b[4]);
    or d5(y[5],a[5],b[5]);
    or d6(y[6],a[6],b[6]);
    or d7(y[7],a[7],b[7]);
    or d8(y[8],a[8],b[8]);
    or d9(y[9],a[9],b[9]);
    or d10(y[10],a[10],b[10]);
    or d11(y[11],a[11],b[11]);
    or d12(y[12],a[12],b[12]);
    or d13(y[13],a[13],b[13]);
    or d14(y[14],a[14],b[14]);
    or d15(y[15],a[15],b[15]);
    or d16(y[16],a[16],b[16]);
    or d17(y[17],a[17],b[17]);
    or d18(y[18],a[18],b[18]);
    or d19(y[19],a[19],b[19]);
    or d20(y[20],a[20],b[20]);
    or d21(y[21],a[21],b[21]);
    or d22(y[22],a[22],b[22]);
    or d23(y[23],a[23],b[23]);
    or d24(y[24],a[24],b[24]);
    or d25(y[25],a[25],b[25]);
    or d26(y[26],a[26],b[26]);
    or d27(y[27],a[27],b[27]);
    or d28(y[28],a[28],b[28]);
    or d29(y[29],a[29],b[29]);
    or d30(y[30],a[30],b[30]);
    or d31(y[31],a[31],b[31]); 
endmodule
    
    

