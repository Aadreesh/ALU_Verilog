module exor
(
    output out,
    input a,b
);

    assign out = a ^ b; 

endmodule