`include "not.v"
module not_all
{
    input [31:0] a,
    output [31:0] out
};
    not c0(y[0],a[0]);
    not c1(y[1],a[1]);
    not c2(y[2],a[2]);
    not c3(y[3],a[3]);
    not c4(y[4],a[4]);
    not c5(y[5],a[5]);
    not c6(y[6],a[6]);
    not c7(y[7],a[7]);
    not c8(y[8],a[8]);
    not c9(y[9],a[9]);
    not c10(y[10],a[10]);
    not c11(y[11],a[11]);
    not c12(y[12],a[12]);
    not c13(y[13],a[13]);
    not c14(y[14],a[14]);
    not c15(y[15],a[15]);
    not c16(y[16],a[16]);
    not c17(y[17],a[17]);
    not c18(y[18],a[18]);
    not c19(y[19],a[19]);
    not c20(y[20],a[20]);
    not c21(y[21],a[21]);
    not c22(y[22],a[22]);
    not c23(y[23],a[23]);
    not c24(y[24],a[24]);
    not c25(y[25],a[25]);
    not c26(y[26],a[26]);
    not c27(y[27],a[27]);
    not c28(y[28],a[28]);
    not c29(y[29],a[29]);
    not c30(y[30],a[30]);
    not c31(y[31],a[31]);
endmodule
    
    

