`include "and.v"
module and_gate4
{
    input [3:0] a, b,
    output [3:0] out
};
    and a0(y[0],a[0],b[0]);
    and a1(y[1],a[1],b[1]);
    and a2(y[2],a[2],b[2);
    and a3(y[3],a[3],b[3]);
endmodule
    
    

