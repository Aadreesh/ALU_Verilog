module not
{
    output out,
    input a ;
};

    assign out = ~a; 

endmodule