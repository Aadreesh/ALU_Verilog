`include "exor.v"
module exor_all
{
    input [31:0] a, b,
    output [31:0] out
};
    exor b0(y[0],a[0],b[0]);
    exor b1(y[1],a[1],b[1]);
    exor b2(y[2],a[2],b[2);
    exor b3(y[3],a[3],b[3]);
    exor b4(y[4],a[4],b[4]);
    exor b5(y[5],a[5],b[5]);
    exor b6(y[6],a[6],b[6]);
    exor b7(y[7],a[7],b[7]);
    exor b8(y[8],a[8],b[8]);
    exor b9(y[9],a[9],b[9]);
    exor b10(y[10],a[10],b[10]);
    exor b11(y[11],a[11],b[11]);
    exor b12(y[12],a[12],b[12]);
    exor b13(y[13],a[13],b[13]);
    exor b14(y[14],a[14],b[14]);
    exor b15(y[15],a[15],b[15]);
    exor b16(y[16],a[16],b[16]);
    exor b17(y[17],a[17],b[17]);
    exor b18(y[18],a[18],b[18]);
    exor b19(y[19],a[19],b[19]);
    exor b20(y[20],a[20],b[20]);
    exor b21(y[21],a[21],b[21]);
    exor b22(y[22],a[22],b[22]);
    exor b23(y[23],a[23],b[23]);
    exor b24(y[24],a[24],b[24]);
    exor b25(y[25],a[25],b[25]);
    exor b26(y[26],a[26],b[26]);
    exor b27(y[27],a[27],b[27]);
    exor b28(y[28],a[28],b[28]);
    exor b29(y[29],a[29],b[29]);
    exor b30(y[30],a[30],b[30]);
    exor b31(y[31],a[31],b[31]);
endmodule
    
    

